module full_adder()