module fourbit_s()